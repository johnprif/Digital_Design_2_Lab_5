library verilog;
use verilog.vl_types.all;
entity full_adder_8_vlg_vec_tst is
end full_adder_8_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity MyLatch_vlg_vec_tst is
end MyLatch_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity REG_8_vlg_vec_tst is
end REG_8_vlg_vec_tst;

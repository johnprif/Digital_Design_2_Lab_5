library verilog;
use verilog.vl_types.all;
entity exercise_B_vlg_vec_tst is
end exercise_B_vlg_vec_tst;
